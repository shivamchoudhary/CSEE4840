library verilog;
use verilog.vl_types.all;
entity SoCKit_Top is
    port(
        AUD_ADCDAT      : in     vl_logic;
        AUD_ADCLRCK     : inout  vl_logic;
        AUD_BCLK        : inout  vl_logic;
        AUD_DACLRCK     : inout  vl_logic;
        AUD_I2C_SDAT    : inout  vl_logic;
        AUD_I2C_SCLK    : out    vl_logic;
        AUD_DACDAT      : out    vl_logic;
        AUD_MUTE        : out    vl_logic;
        AUD_XCK         : out    vl_logic;
        FAN_CTRL        : out    vl_logic;
        HSMC_CLKIN_n    : in     vl_logic_vector(2 downto 1);
        HSMC_CLKIN_p    : in     vl_logic_vector(2 downto 1);
        HSMC_CLKOUT_n   : out    vl_logic_vector(2 downto 1);
        HSMC_CLKOUT_p   : out    vl_logic_vector(2 downto 1);
        HSMC_CLK_IN0    : in     vl_logic;
        HSMC_CLK_OUT0   : out    vl_logic;
        HSMC_D          : inout  vl_logic_vector(3 downto 0);
        HSMC_RX_n       : inout  vl_logic_vector(16 downto 0);
        HSMC_RX_p       : inout  vl_logic_vector(16 downto 0);
        HSMC_TX_n       : inout  vl_logic_vector(16 downto 0);
        HSMC_TX_p       : inout  vl_logic_vector(16 downto 0);
        HSMC_SDA        : inout  vl_logic;
        HSMC_SCL        : out    vl_logic;
        IRDA_RXD        : in     vl_logic;
        KEY             : in     vl_logic_vector(3 downto 0);
        LED             : out    vl_logic_vector(3 downto 0);
        OSC_50_B3B      : in     vl_logic;
        OSC_50_B4A      : in     vl_logic;
        OSC_50_B5B      : in     vl_logic;
        OSC_50_B8A      : in     vl_logic;
        PCIE_PERST_n    : in     vl_logic;
        PCIE_WAKE_n     : in     vl_logic;
        RESET_n         : in     vl_logic;
        SI5338_SCL      : inout  vl_logic;
        SI5338_SDA      : inout  vl_logic;
        SW              : in     vl_logic_vector(3 downto 0);
        TEMP_CS_n       : out    vl_logic;
        TEMP_DIN        : out    vl_logic;
        TEMP_SCLK       : out    vl_logic;
        TEMP_DOUT       : in     vl_logic;
        USB_B2_CLK      : in     vl_logic;
        USB_OE_n        : in     vl_logic;
        USB_RD_n        : in     vl_logic;
        USB_WR_n        : in     vl_logic;
        USB_RESET_n     : in     vl_logic;
        USB_B2_DATA     : inout  vl_logic_vector(7 downto 0);
        USB_EMPTY       : out    vl_logic;
        USB_FULL        : out    vl_logic;
        USB_SCL         : inout  vl_logic;
        USB_SDA         : inout  vl_logic;
        VGA_R           : out    vl_logic_vector(7 downto 0);
        VGA_G           : out    vl_logic_vector(7 downto 0);
        VGA_B           : out    vl_logic_vector(7 downto 0);
        VGA_CLK         : out    vl_logic;
        VGA_HS          : out    vl_logic;
        VGA_VS          : out    vl_logic;
        VGA_BLANK_n     : out    vl_logic;
        VGA_SYNC_n      : out    vl_logic
    );
end SoCKit_Top;
